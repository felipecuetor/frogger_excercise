//=======================================================
//  MODULE Definition
//=======================================================
module REGDI_NV#(parameter NV_1_REG, 	parameter NV_2_REG, 	parameter NV_3_REG, 	parameter NV_4_REG ) 
(
//////////// OUTPUTS //////////
   REGDI_NV_DATAPARALLEL_OUT,
//////////// INPUTS //////////
	REGDI_NV_CLOCK,
	REGDI_NV_RESET,
	REGDI_NV_NVL_IN,
	REGDI_NV_CN_IN
);
//=======================================================
//  PARAMETER declarations
//=======================================================
	parameter DATAWIDTH_BUS = 8;
	parameter CLOCK0_DATAWITH= 3; //RAPIDO
	parameter CLOCK1_DATAWITH= 4; //NORMAL
	parameter CLOCK2_DATAWITH= 5; //LENTO
	parameter DATAWIDTH_SELECTOR=2;
	parameter DATAWIDTH_NIVEL=2;
//=======================================================
//  PORT declarations
//=======================================================
	output [DATAWIDTH_BUS-1:0] REGDI_NV_DATAPARALLEL_OUT;
	input	REGDI_NV_CLOCK;
	input REGDI_NV_RESET;
	input [DATAWIDTH_NIVEL-1:0] REGDI_NV_NVL_IN;
	input REGDI_NV_CN_IN;
//=======================================================
//  REG/WIRE declarations
//=======================================================
	wire REGDI_NV_LOAD;
	wire REGDI_NV_SHIFT;
	wire REGDI_NV_LOADED;
	wire [DATAWIDTH_BUS-1:0] REGDI_NV_DATAPARALLEL_BUS;
	
	wire REGDI_NV_RECLOCK0;
	wire REGDI_NV_RECLOCK1;
	wire REGDI_NV_RECLOCK2;
	wire [DATAWIDTH_SELECTOR-1:0] REGDI_NV_CLOCK_SELECT;
	wire REGDI_NV_CLOCK_SELECTED;
	wire REGDI_NV_RECLOCK0_HAB;
	wire REGDI_NV_RECLOCK1_HAB;
	wire REGDI_NV_RECLOCK2_HAB;
	
//=======================================================
//  Structural coding
//=======================================================
	
	SC_REGDI #(.DATAWIDTH_BUS(DATAWIDTH_BUS)) 
	SC_REGDI_u0 (
// port map - connection between master ports and signals/registers   
	.SC_REGDI_DATAPARALLEL_BUS_OUT(REGDI_NV_DATAPARALLEL_OUT),
	.SC_REGDI_CLOCK(REGDI_NV_CLOCK_SELECTED),
	.SC_REGDI_RESET(REGDI_NV_RESET),
	.SC_REGDI_DATAPARALLEL_BUS_IN(REGDI_NV_DATAPARALLEL_BUS),
	.SC_REGDI_LOAD(REGDI_NV_LOAD),
	.SC_REGDI_LOADED(REGDI_NV_LOADED),
	.SC_REGDI_SHIFT(REGDI_NV_SHIFT)
);

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK0_DATAWITH))
	SC_RECLOCK_u0(
	.SC_RECLOCK_Out(REGDI_NV_RECLOCK0),
	.SC_RECLOCK_CLOCK_50(REGDI_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDI_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDI_NV_RECLOCK0_HAB)
);	

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK1_DATAWITH))
	SC_RECLOCK_u1(
	.SC_RECLOCK_Out(REGDI_NV_RECLOCK1),
	.SC_RECLOCK_CLOCK_50(REGDI_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDI_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDI_NV_RECLOCK1_HAB)
);

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK2_DATAWITH))
	SC_RECLOCK_u2(
	.SC_RECLOCK_Out(REGDI_NV_RECLOCK2),
	.SC_RECLOCK_CLOCK_50(REGDI_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDI_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDI_NV_RECLOCK2_HAB)
);


MUXX41 #(.DATAWIDTH_SELECTOR(DATAWIDTH_SELECTOR))
 MUXX41_u0(
	.MUXX41_Z_BIT_OUT(REGDI_NV_CLOCK_SELECTED),
	.MUXX41_SELECT_BUS_IN(REGDI_NV_CLOCK_SELECT),
	.MUXX41_IN0(REGDI_NV_CLOCK),
	.MUXX41_IN1(REGDI_NV_RECLOCK2),
	.MUXX41_IN2(REGDI_NV_RECLOCK1),
	.MUXX41_IN3(REGDI_NV_RECLOCK0)
);	
	SC_STATEMACHINE_NVE #(.DATAWIDTH_BUS(DATAWIDTH_BUS), .NV_1_REG(NV_1_REG), .NV_2_REG(NV_2_REG), .NV_3_REG(NV_3_REG), .NV_4_REG(NV_4_REG))
	SC_STATEMACHINE_NVE_u0(
	.SC_STATEMACHINE_NVE_LOAD_OUT(REGDI_NV_LOAD),
	.SC_STATEMACHINE_NVE_SHIFT_OUT(REGDI_NV_SHIFT),
	.SC_STATEMACHINE_NVE_HAB_CLOCK0_OUT(REGDI_NV_RECLOCK0_HAB),
	.SC_STATEMACHINE_NVE_HAB_CLOCK1_OUT(REGDI_NV_RECLOCK1_HAB),
	.SC_STATEMACHINE_NVE_HAB_CLOCK2_OUT(REGDI_NV_RECLOCK2_HAB),
	.SC_STATEMACHINE_NVE_CLOCK_SELECT(REGDI_NV_CLOCK_SELECT),
	.SC_STATEMACHINE_NVE_REGNIVEL_OUT(REGDI_NV_DATAPARALLEL_BUS),
	.SC_STATEMACHINE_NVE_NVL_IN(REGDI_NV_NVL_IN),
	.SC_STATEMACHINE_NVE_CN_IN(REGDI_NV_CN_IN),
	.SC_STATEMACHINE_NVE_LOADED_IN(REGDI_NV_LOADED),
	.SC_STATEMACHINE_NVE_CLOCK_50(REGDI_NV_CLOCK),
	.SC_STATEMACHINE_NVE_RESET(REGDI_NV_RESET)
);	
  
endmodule

