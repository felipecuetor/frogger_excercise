//=======================================================
//  MODULE Definition
//=======================================================
module JUEGO (
//////////// OUTPUTS //////////
   JUEGO_7_OUT,
   JUEGO_6_OUT,
	JUEGO_5_OUT,
	JUEGO_4_OUT,
	JUEGO_3_OUT,
	JUEGO_2_OUT,
	JUEGO_1_OUT,
	JUEGO_0_OUT, 
//////////// INPUTS //////////
	JUEGO_CLOCK,
	JUEGO_RESET,	
	JUEGO_START,
	JUEGO_LEFT,
	JUEGO_RIGHT,
	JUEGO_UP,
	JUEGO_DOWN
	
);
//=======================================================
//  PARAMETER declarations
//=======================================================
		parameter DATAWIDTH_BUS = 8;
		parameter DATAWIDTH_ESTADO = 3;
		parameter DATAWIDTH_POS = 3;
		parameter DATAWIDTH_NV = 2;
//=======================================================
//  PORT declarations
//=======================================================
	output wire[DATAWIDTH_BUS-1:0] JUEGO_7_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_6_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_5_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_4_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_3_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_2_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_1_OUT;
	output wire[DATAWIDTH_BUS-1:0] JUEGO_0_OUT;
	input wire JUEGO_CLOCK;
	input wire JUEGO_RESET;	
	input wire JUEGO_START;
	input wire JUEGO_LEFT;
	input wire JUEGO_RIGHT;
	input wire JUEGO_UP;
	input wire JUEGO_DOWN;
	
//=======================================================
//  REG/WIRE declarations
//=======================================================		

	wire [DATAWIDTH_BUS-1:0] JUEGONV_7;
	
	wire [DATAWIDTH_BUS-1:0] JUEGONV_6;
	wire [DATAWIDTH_BUS-1:0] JUEGONV_5;
	wire [DATAWIDTH_BUS-1:0] JUEGONV_4;
	wire [DATAWIDTH_BUS-1:0] JUEGONV_3;
	wire [DATAWIDTH_BUS-1:0] JUEGONV_2;
	wire [DATAWIDTH_BUS-1:0] JUEGONV_1;
	
	wire [DATAWIDTH_BUS-1:0] JDATA_7;
	wire [DATAWIDTH_BUS-1:0] JDATA_6;
	wire [DATAWIDTH_BUS-1:0] JDATA_5;
	wire [DATAWIDTH_BUS-1:0] JDATA_4;
	wire [DATAWIDTH_BUS-1:0] JDATA_3;
	wire [DATAWIDTH_BUS-1:0] JDATA_2;
	wire [DATAWIDTH_BUS-1:0] JDATA_1;
	wire [DATAWIDTH_BUS-1:0] JDATA_0;
	
	
	wire [DATAWIDTH_NV-1:0] JUEGO_W_NVL;
	wire JUEGO_W_CN;
	wire [DATAWIDTH_ESTADO-1:0] JUEGO_W_ESTADO;
   wire [DATAWIDTH_POS-1:0] JUEGO_W_POSX;
	wire [DATAWIDTH_POS-1:0] JUEGO_W_POSY;
	wire JUEGO_W_PERDIO;
	wire JUEGO_W_GANO;
	wire JUEGO_RANAINI;
		
//=======================================================
//  Structural coding
//=======================================================
	MENU_PRINCIPAL
	MENU_PRINCIPAL_u0 (
	.MP_ESTADO_OUT(JUEGO_W_ESTADO),
	.MP_NVL_OUT(JUEGO_W_NVL),
	.MP_CN_OUT(JUEGO_W_CN),
	.MP_GANO(JUEGO_W_GANO),
	.MP_PERDIO(JUEGO_W_PERDIO),
	.MP_DOWN(JUEGO_DOWN),
	.MP_UP(JUEGO_UP),
	.MP_START(JUEGO_START),
	.MP_CLOCK_50(JUEGO_CLOCK),
	.MP_RESET(JUEGO_RESET)
	);
	
	NIVEL_VEHICULOS
	NIVEL_VEHICULOS_u0 (
	.NVE_REG_5_OUT(JUEGONV_6),
	.NVE_REG_4_OUT(JUEGONV_5),
	.NVE_REG_3_OUT(JUEGONV_4),
	.NVE_REG_2_OUT(JUEGONV_3),
	.NVE_REG_1_OUT(JUEGONV_2),
	.NVE_REG_0_OUT(JUEGONV_1),
	.NVE_CLOCK(JUEGO_CLOCK),
	.NVE_RESET(JUEGO_RESET),
	.NVE_ESTADO_IN(JUEGO_W_ESTADO),
	.NVE_NV_IN(JUEGO_W_NVL),
	.NVE_CN_IN(JUEGO_W_CN)
	); 
	
	CONTROL_RANAS
	CONTROL_RANAS_u0(
	.CR_GANO_JC_OUT(JUEGO_W_GANO),
	.CR_RANA_INI_OUT(JUEGO_RANAINI),
	.CR_POSY_IN(JUEGO_W_POSY),
	.CR_PERDIO_IN(JUEGO_W_PERDIO),
	.CR_ESTADO_IN(JUEGO_W_ESTADO),
	.CR_CLOCK_50(JUEGO_CLOCK),
	.CR_RESET(JUEGO_RESET)
	);
	
	CONTROL_CASAS
	CONTROL_CASAS_u0(
	.CC_REG7_OUT(JUEGONV_7),
	.CC_POSX_IN(JUEGO_W_POSX),
	.CC_POSY_IN(JUEGO_W_POSY),
	.CC_PERDIO_IN(JUEGO_W_PERDIO),
	.CC_ESTADO_IN(JUEGO_W_ESTADO),
	.CC_CLOCK_50(JUEGO_CLOCK),
	.CC_RESET(JUEGO_RESET)
	);
	
	COLISION
	COLISION_u0 (
	.CO_PERDIO_OUT(JUEGO_W_PERDIO),
	.CO_POSX_IN(JUEGO_W_POSX),
	.CO_POSY_IN(JUEGO_W_POSY),
	.CO_VEH7_IN(JUEGONV_7),
	.CO_VEH6_IN(JUEGONV_6),
	.CO_VEH5_IN(JUEGONV_5),
	.CO_VEH4_IN(JUEGONV_4),
	.CO_VEH3_IN(JUEGONV_3),
	.CO_VEH2_IN(JUEGONV_2),
	.CO_VEH1_IN(JUEGONV_1)
);

	RANA 
	RANA_u0(
    .RANA_7_OUT(JDATA_7),
	 .RANA_6_OUT(JDATA_6),
	 .RANA_5_OUT(JDATA_5),
	 .RANA_4_OUT(JDATA_4),
	 .RANA_3_OUT(JDATA_3),
	 .RANA_2_OUT(JDATA_2),
	 .RANA_1_OUT(JDATA_1),
	 .RANA_0_OUT(JDATA_0),
	 .PXRANA_OUT(JUEGO_W_POSX),
	 .PYRANA_OUT(JUEGO_W_POSY),
	 .RANA_CLOCK(JUEGO_CLOCK),
	 .RANA_RESET(JUEGO_RESET),
	 .RANA_INI(JUEGO_RANAINI),
	 .RANA_LEFT(JUEGO_LEFT),
	 .RANA_RIGHT(JUEGO_RIGHT),
	 .RANA_UP(JUEGO_UP),
	 .RANA_DOWN(JUEGO_DOWN),
	 .VEH7_IN(JUEGONV_7),
	 .VEH6_IN(JUEGONV_6),
	 .VEH5_IN(JUEGONV_5),
	 .VEH4_IN(JUEGONV_4),
	 .VEH3_IN(JUEGONV_3),
	 .VEH2_IN(JUEGONV_2),
	 .VEH1_IN(JUEGONV_1)
	);
	
	PINTAR_MATRIZ 
	PINTAR_MATRIZ_u0 (
	.PINTAR_7_OUT(JUEGO_7_OUT),
	.PINTAR_6_OUT(JUEGO_6_OUT),
	.PINTAR_5_OUT(JUEGO_5_OUT),
	.PINTAR_4_OUT(JUEGO_4_OUT),
	.PINTAR_3_OUT(JUEGO_3_OUT),
	.PINTAR_2_OUT(JUEGO_2_OUT),
	.PINTAR_1_OUT(JUEGO_1_OUT),
	.PINTAR_0_OUT(JUEGO_0_OUT),
	.PINTAR_J7_IN(JDATA_7),
	.PINTAR_J6_IN(JDATA_6),
	.PINTAR_J5_IN(JDATA_5),
	.PINTAR_J4_IN(JDATA_4),
	.PINTAR_J3_IN(JDATA_3),
	.PINTAR_J2_IN(JDATA_2),
	.PINTAR_J1_IN(JDATA_1),
	.PINTAR_J0_IN(JDATA_0),
	.PINTAR_MENU_PRINCIPAL_ESTADO_IN(JUEGO_W_ESTADO)
);
	
										
endmodule 