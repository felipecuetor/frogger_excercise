//=======================================================
//  MODULE Definition
//=======================================================
module REG_NV
(
//////////// OUTPUTS //////////
   REGDD_NV_DATAPARALLEL_OUT,
	REGDI_NV_DATAPARALLEL_OUT,
//////////// INPUTS //////////
	REG_NV_CLOCK,
	REG_NV_RESET,
	REG_NV_NVL_IN,
	REG_NV_CN_IN
);
//=======================================================
//  PARAMETER declarations
//=======================================================
	//VELOCIDADES
	parameter VEL0_DATAWITH= 3; //RAPIDO
	parameter VEL1_DATAWITH= 4; //NORMAL
	parameter VEL2_DATAWITH= 5; //LENTO
	//NIVELES
	parameter NV_1_REGD =   8'b11000000;
	parameter NV_2_REGD =	8'b11100000;
	parameter NV_3_REGD =	8'b11110000;
	parameter NV_4_REGD =	8'b11111000;
	parameter NV_1_REGI =	8'b00000000;
	parameter NV_2_REGI =	8'b00000011;
	parameter NV_3_REGI =	8'b00000111;
	parameter NV_4_REGI =	8'b00001111;
	parameter DATAWIDTH_BUS = 8;
	parameter DATAWIDTH_SELECTOR=2;
	parameter DATAWIDTH_NVL=2;
//=======================================================
//  PORT declarations
//=======================================================
	output [DATAWIDTH_BUS-1:0] REGDD_NV_DATAPARALLEL_OUT;
	output [DATAWIDTH_BUS-1:0] REGDI_NV_DATAPARALLEL_OUT;
	input	REG_NV_CLOCK;
	input REG_NV_RESET;
	input [DATAWIDTH_NVL-1:0] REG_NV_NVL_IN;
	input REG_NV_CN_IN;
//=======================================================
//  REG/WIRE declarations
//=======================================================
	wire REG_NV_LOAD_SHIFT;
	wire [DATAWIDTH_BUS-1:0] REGDD_NV_DATAPARALLEL_BUS;
	wire [DATAWIDTH_BUS-1:0] REGDI_NV_DATAPARALLEL_BUS;
	wire REG_NV_VEL0;
	wire REG_NV_VEL1;
	wire REG_NV_VEL2;
	wire [DATAWIDTH_SELECTOR-1:0] REG_NV_VEL_SELECT;
	wire REG_NV_VEL_SELECTED;
	wire REG_NV_VEL0_HAB;
	wire REG_NV_VEL1_HAB;
	wire REG_NV_VEL2_HAB;
	
//=======================================================
//  Structural coding
//=======================================================

	SC_REGDI #(.DATAWIDTH_BUS(DATAWIDTH_BUS)) 
	SC_REGDI_u0 (  
	.SC_REGDI_DATAPARALLEL_BUS_OUT(REGDI_NV_DATAPARALLEL_OUT),
	.SC_REGDI_CLOCK(REG_NV_CLOCK),
	.SC_REGDI_RESET(REG_NV_RESET),
	.SC_REGDI_VEL(REG_NV_VEL_SELECTED),
	.SC_REGDI_LOAD_SHIFT(REG_NV_LOAD_SHIFT),
	.SC_REGDI_DATAPARALLEL_BUS_IN(REGDI_NV_DATAPARALLEL_BUS)
);
	
	SC_REGDD #(.DATAWIDTH_BUS(DATAWIDTH_BUS)) 
	SC_REGDD_u0 (
	.SC_REGDD_DATAPARALLEL_BUS_OUT(REGDD_NV_DATAPARALLEL_OUT),
	.SC_REGDD_CLOCK(REG_NV_CLOCK),
	.SC_REGDD_RESET(REG_NV_RESET),
	.SC_REGDD_VEL(REG_NV_VEL_SELECTED),
	.SC_REGDD_LOAD_SHIFT(REG_NV_LOAD_SHIFT),
	.SC_REGDD_DATAPARALLEL_BUS_IN(REGDD_NV_DATAPARALLEL_BUS)
);



	SC_VEL #(.VEL_DATAWITH(VEL0_DATAWITH))
	SC_VEL_u0(
	.SC_VEL_OUT(REG_NV_VEL0),
	.SC_VEL_CLOCK_50(REG_NV_CLOCK),
	.SC_VEL_RESET(REG_NV_RESET),
	.SC_VEL_HAB_IN(REG_NV_VEL0_HAB)
);	

	SC_VEL #(.VEL_DATAWITH(VEL1_DATAWITH))
	SC_VEL_u1(
	.SC_VEL_OUT(REG_NV_VEL1),
	.SC_VEL_CLOCK_50(REG_NV_CLOCK),
	.SC_VEL_RESET(REG_NV_RESET),
	.SC_VEL_HAB_IN(REG_NV_VEL1_HAB)
);

	SC_VEL #(.VEL_DATAWITH(VEL2_DATAWITH))
	SC_VEL_u2(
	.SC_VEL_OUT(REG_NV_VEL2),
	.SC_VEL_CLOCK_50(REG_NV_CLOCK),
	.SC_VEL_RESET(REG_NV_RESET),
	.SC_VEL_HAB_IN(REG_NV_VEL2_HAB)
);


MUXX41 #(.DATAWIDTH_SELECTOR(DATAWIDTH_SELECTOR))
 MUXX41_u0(
	.MUXX41_Z_BIT_OUT(REG_NV_VEL_SELECTED),
	.MUXX41_SELECT_BUS_IN(REG_NV_VEL_SELECT),
	.MUXX41_IN0(1'b0),
	.MUXX41_IN1(REG_NV_VEL2),
	.MUXX41_IN2(REG_NV_VEL1),
	.MUXX41_IN3(REG_NV_VEL0)
);	
	SC_STATEMACHINE_NVE #(.DATAWIDTH_BUS(DATAWIDTH_BUS), .NV_1_REGD(NV_1_REGD), .NV_2_REGD(NV_2_REGD), .NV_3_REGD(NV_3_REGD), .NV_4_REGD(NV_4_REGD), .NV_1_REGI(NV_1_REGI), .NV_2_REGI(NV_2_REGI), .NV_3_REGI(NV_3_REGI), .NV_4_REGI(NV_4_REGI))
	SC_STATEMACHINE_NVE_u0(
	.SC_STATEMACHINE_NVE_LOAD_SHIFT_OUT(REG_NV_LOAD_SHIFT),
	.SC_STATEMACHINE_NVE_VEL_SELECT(REG_NV_VEL_SELECT),
	.SC_STATEMACHINE_NVE_HAB_VEL0_OUT(REG_NV_VEL0_HAB),
	.SC_STATEMACHINE_NVE_HAB_VEL1_OUT(REG_NV_VEL1_HAB),
	.SC_STATEMACHINE_NVE_HAB_VEL2_OUT(REG_NV_VEL2_HAB),
	.SC_STATEMACHINE_NVE_REGDNIVEL_OUT(REGDD_NV_DATAPARALLEL_BUS),
	.SC_STATEMACHINE_NVE_REGINIVEL_OUT(REGDI_NV_DATAPARALLEL_BUS),
	.SC_STATEMACHINE_NVE_NVL_IN(REG_NV_NVL_IN),
	.SC_STATEMACHINE_NVE_CN_IN(REG_NV_CN_IN),
	.SC_STATEMACHINE_NVE_CLOCK_50(REG_NV_CLOCK),
	.SC_STATEMACHINE_NVE_RESET(REG_NV_RESET)
);	
  
endmodule

