//=======================================================
//  MODULE Definition
//=======================================================
module REGDD_NV#(parameter NV_1_REG, 	parameter NV_2_REG, 	parameter NV_3_REG, 	parameter NV_4_REG ) 
(
//////////// OUTPUTS //////////
   REGDD_NV_DATAPARALLEL_OUT,
//////////// INPUTS //////////
	REGDD_NV_CLOCK,
	REGDD_NV_RESET,
	REGDD_NV_NVL_IN,
	REGDD_NV_CN_IN
);
//=======================================================
//  PARAMETER declarations
//=======================================================
	parameter DATAWIDTH_BUS = 8;
	parameter CLOCK0_DATAWITH= 3; //RAPIDO
	parameter CLOCK1_DATAWITH= 4; //NORMAL
	parameter CLOCK2_DATAWITH= 5; //LENTO
	parameter DATAWIDTH_SELECTOR=2;
	parameter DATAWIDTH_NVL=2;
//=======================================================
//  PORT declarations
//=======================================================
	output [DATAWIDTH_BUS-1:0] REGDD_NV_DATAPARALLEL_OUT;
	input	REGDD_NV_CLOCK;
	input REGDD_NV_RESET;
	input [DATAWIDTH_NVL-1:0] REGDD_NV_NVL_IN;
	input REGDD_NV_CN_IN;
//=======================================================
//  REG/WIRE declarations
//=======================================================
	wire REGDD_NV_LOAD;
	wire REGDD_NV_SHIFT;
	wire REGDD_NV_LOADED;
	wire [DATAWIDTH_BUS-1:0] REGDD_NV_DATAPARALLEL_BUS;
	
	wire REGDD_NV_RECLOCK0;
	wire REGDD_NV_RECLOCK1;
	wire REGDD_NV_RECLOCK2;
	wire [DATAWIDTH_SELECTOR-1:0] REGDD_NV_CLOCK_SELECT;
	wire REGDD_NV_CLOCK_SELECTED;
	wire REGDD_NV_RECLOCK0_HAB;
	wire REGDD_NV_RECLOCK1_HAB;
	wire REGDD_NV_RECLOCK2_HAB;
	
//=======================================================
//  Structural coding
//=======================================================
	
	SC_REGDD #(.DATAWIDTH_BUS(DATAWIDTH_BUS)) 
	SC_REGDD_u0 (
// port map - connection between master ports and signals/registers   
	.SC_REGDD_DATAPARALLEL_BUS_OUT(REGDD_NV_DATAPARALLEL_OUT),
	.SC_REGDD_CLOCK(REGDD_NV_CLOCK_SELECTED),
	.SC_REGDD_RESET(REGDD_NV_RESET),
	.SC_REGDD_DATAPARALLEL_BUS_IN(REGDD_NV_DATAPARALLEL_BUS),
	.SC_REGDD_LOAD(REGDD_NV_LOAD),
	.SC_REGDD_LOADED(REGDD_NV_LOADED),
	.SC_REGDD_SHIFT(REGDD_NV_SHIFT)
);

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK0_DATAWITH))
	SC_RECLOCK_u0(
	.SC_RECLOCK_Out(REGDD_NV_RECLOCK0),
	.SC_RECLOCK_CLOCK_50(REGDD_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDD_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDD_NV_RECLOCK0_HAB)
);	

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK1_DATAWITH))
	SC_RECLOCK_u1(
	.SC_RECLOCK_Out(REGDD_NV_RECLOCK1),
	.SC_RECLOCK_CLOCK_50(REGDD_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDD_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDD_NV_RECLOCK1_HAB)
);

	SC_RECLOCK #(.CLOCK_DATAWITH(CLOCK2_DATAWITH))
	SC_RECLOCK_u2(
	.SC_RECLOCK_Out(REGDD_NV_RECLOCK2),
	.SC_RECLOCK_CLOCK_50(REGDD_NV_CLOCK),
	.SC_RECLOCK_RESET(REGDD_NV_RESET),
	.SC_RECLOCK_HAB_IN(REGDD_NV_RECLOCK2_HAB)
);


MUXX41 #(.DATAWIDTH_SELECTOR(DATAWIDTH_SELECTOR))
 MUXX41_u0(
	.MUXX41_Z_BIT_OUT(REGDD_NV_CLOCK_SELECTED),
	.MUXX41_SELECT_BUS_IN(REGDD_NV_CLOCK_SELECT),
	.MUXX41_IN0(REGDD_NV_CLOCK),
	.MUXX41_IN1(REGDD_NV_RECLOCK2),
	.MUXX41_IN2(REGDD_NV_RECLOCK1),
	.MUXX41_IN3(REGDD_NV_RECLOCK0)
);	
	SC_STATEMACHINE_NVE #(.DATAWIDTH_BUS(DATAWIDTH_BUS), .NV_1_REG(NV_1_REG), .NV_2_REG(NV_2_REG), .NV_3_REG(NV_3_REG), .NV_4_REG(NV_4_REG))
	SC_STATEMACHINE_NVE_u0(
	.SC_STATEMACHINE_NVE_LOAD_OUT(REGDD_NV_LOAD),
	.SC_STATEMACHINE_NVE_SHIFT_OUT(REGDD_NV_SHIFT),
	.SC_STATEMACHINE_NVE_HAB_CLOCK0_OUT(REGDD_NV_RECLOCK0_HAB),
	.SC_STATEMACHINE_NVE_HAB_CLOCK1_OUT(REGDD_NV_RECLOCK1_HAB),
	.SC_STATEMACHINE_NVE_HAB_CLOCK2_OUT(REGDD_NV_RECLOCK2_HAB),
	.SC_STATEMACHINE_NVE_CLOCK_SELECT(REGDD_NV_CLOCK_SELECT),
	.SC_STATEMACHINE_NVE_REGNIVEL_OUT(REGDD_NV_DATAPARALLEL_BUS),
	.SC_STATEMACHINE_NVE_NVL_IN(REGDD_NV_NVL_IN),
	.SC_STATEMACHINE_NVE_CN_IN(REGDD_NV_CN_IN),
	.SC_STATEMACHINE_NVE_LOADED_IN(REGDD_NV_LOADED),
	.SC_STATEMACHINE_NVE_CLOCK_50(REGDD_NV_CLOCK),
	.SC_STATEMACHINE_NVE_RESET(REGDD_NV_RESET)
);	
  
endmodule

